\m5_TLV_version 1d: tl-x.org
\m5


   //use(m5-1.0)   /// uncomment to use M5 macro library.
\SV
   
   m5_makerchip_module   // (Expanded in Nav-TLV pane.)

\TLV
   $reset = *reset;

    $sum[31:0] = $val1[31:0] + $val2[31:0];
    $diff[31:0] = $val1[31:0] - $val2[31:0];
    $prod[31:0] = $val1[31:0] * $val2[31:0];
    $quot[31:0] = $val1[31:0] / $val2[31:0];
    $out[31:0] = $op[0] ? $sum : $op[1] ? $diff : $op[2] ? $prod : $qout ;

   // Assert these to end simulation (before the cycle limit).
   *passed = *cyc_cnt > 40;
   *failed = 1'b0;
\SV
   endmodule
